module student_circuit_Q1 (
          input clk, clear,
          input [7:0] cct_input,
          output reg [7:0] cct_output
			 );


endmodule
