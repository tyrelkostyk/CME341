module student_circuit_Q3b (
          input clk, clear,
          input [7:0] cct_input,
          output reg [7:0] cct_output
			 );



endmodule
