module student_circuit (
          input clk, clear,
          input [7:0] cct_input,
          output [7:0] cct_output  // for the answers
			 );


// student_circuit_Q1 the_cct(			 
// student_circuit_Q2 the_cct(			 
// student_circuit_Q3A the_cct(	
// student_circuit_Q3B the_cct(		 
// student_circuit_Q4 the_cct(	
 student_circuit_Q5 the_cct(			 
          .clk(clk), .clear(clear),
          .cct_input(cct_input),
          .cct_output(cct_output) );
  
  
endmodule